maton@Ubuntu22.6133:1770404027