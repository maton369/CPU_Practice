-- fetch.vhd（詳細コメント版：命令フェッチ段 / PROM（命令ROM）読み出し）
--
-- 【このモジュールの目的（CPU設計観点）】
-- - CPUの Fetch 段として、プログラムカウンタ PC（ここでは P_COUNT）を使い、
--   命令ROM（PROM）から命令ワードを読み出して `PROM_OUT` に出力する。
-- - 自作CPUにおけるフェッチ段は、以下の2点を満たす必要がある：
--   1) PCが指す命令を確実に取り出す（アドレス→命令の対応）
--   2) 取り出した命令を “次段（Decode）で安定して読めるタイミング” で提示する
--
-- 【設計上の特徴（この教材CPUの事情）】
-- - PROMは「配列 + constant 初期化」で実装されており、RAMではなくROM相当である。
-- - 命令語は 15bit 固定（std_logic_vector(14 downto 0)）。
-- - アドレス空間は 0〜15（16語）だけを使う簡易PROMで、
--   PCの下位4bit（P_COUNT(3 downto 0)）で参照している。
--   つまり、このCPUは実験用に “16命令だけ入る小さいプログラム” を実行する構成である。
--
-- 【フェッチ段のアルゴリズム（1サイクル動作）】
-- - CLK_FT（Fetch用ステージクロック）の立ち上がりで、
--   PROM[ PC ] を読み出し PROM_OUT にラッチする。
-- - これにより、次のDecode段（CLK_DC）では PROM_OUT が安定した入力として扱える。
--
-- 【注意：P_COUNT(3 downto 0) を使う意味】
-- - MEM の配列サイズが 16 (=2^4) なので、アドレスとして 4bit しか使っていない。
-- - 上位ビット P_COUNT(7 downto 4) はこのfetchでは無視される。
--   そのため、PCが16以上になってもアドレスは下位4bitで折り返す（モジュロ16動作）になる。
-- - 自作CPUの拡張では、MEMORY を 256語などに拡張し、
--   P_COUNT(7 downto 0) 全体で参照するのが自然になる。
--
-- 【命令ROMの中身（このプログラムが何をするか）】
-- - コメントにある通り、1+2+...+10 の総和（55）を計算し、メモリ(64番地)へ store して停止する。
-- - これは “命令フェッチ→デコード→演算→分岐→ストア→停止” を一通り通るため、
--   CPU bring-up（最初にCPUを動かす試験）用の典型的なスモークテストプログラムになっている。
--
-- 【命令列の流れ（概念）】
--  0: REG0 = 0
--  1: REG1 = 1
--  2: REG2 = 0   （累積値 or 作業レジスタ）
--  3: REG3 = 10  （比較用：上限）
--  8: REG2 = REG2 + REG1   （1ずつ増える値を作る/または加算の一部）
--  9: REG0 = REG0 + REG2   （総和をREG0へ蓄積）
-- 10: MEM[64] = REG0       （結果をI/O相当へ出す想定）
-- 11: if REG2 == REG3 then goto 14
-- 13: goto 8
-- 14: halt
--
-- ここで重要なのは「Fetchが正しく動くと、この“制御フロー”が成立する」という点である。
-- 分岐命令（je/jmp）でPCが変化しても、正しい番地の命令が出てくる必要がある。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- ============================================================
-- entity: Fetch段の外部インタフェース
-- ============================================================
entity fetch is
    port
    (
        -- Fetch段用ステージクロック（clk_genが生成）
        -- この立ち上がりで命令を読み出す。
        CLK_FT   : in  std_logic;

        -- プログラムカウンタ（PC）
        -- exec段で更新され、ここでPROMのアドレスとして使われる。
        P_COUNT  : in  std_logic_vector(7 downto 0);

        -- 命令ROM（PROM）から読み出した命令ワード（15bit）
        -- 次段（decode）へ渡す。
        PROM_OUT : out std_logic_vector(14 downto 0)
    );
end fetch;

-- ============================================================
-- architecture RTL: PROM（命令ROM）を配列で表現し読み出す
-- ============================================================
architecture RTL of fetch is

    -- --------------------------------------------------------
    -- 命令語の型（15bit固定長）
    -- --------------------------------------------------------
    subtype WORD is std_logic_vector(14 downto 0);

    -- --------------------------------------------------------
    -- PROMメモリ型：16語の命令ROM
    -- --------------------------------------------------------
    -- 0〜15 の16エントリだけ持つ超小型PROM。
    type MEMORY is array (0 to 15) of WORD;

    -- --------------------------------------------------------
    -- PROMの中身：固定プログラム
    -- --------------------------------------------------------
    -- CPU動作確認用のプログラム（1+2+...+10=55 の計算＋store＋halt）。
    -- 末尾に nop 相当（全0）も入れている。
    constant MEM : MEMORY :=
        (
            "100100000000000",  -- 0: ldh Reg0, 0   （Reg0の上位8bitへ0をロード）
            "100000000000000",  -- 1: ldl Reg0, 0   （Reg0の下位8bitへ0をロード）=> Reg0=0
            "100100100000000",  -- 2: ldh Reg1, 0
            "100000100000001",  -- 3: ldl Reg1, 1   => Reg1=1
            "100101000000000",  -- 4: ldh Reg2, 0
            "100001000000000",  -- 5: ldl Reg2, 0   => Reg2=0
            "100101100000000",  -- 6: ldh Reg3, 0
            "100001100001010",  -- 7: ldl Reg3, 10  => Reg3=10
            "000101000100000",  -- 8: add Reg2, Reg1 （Reg2 = Reg2 + Reg1）
            "000100001000000",  -- 9: add Reg0, Reg2 （Reg0 = Reg0 + Reg2）=> 総和蓄積
            "111000001000000",  --10: st  Reg0, 64   （結果をRAM/I/Oの64番地へ保存）
            "101001001100000",  --11: cmp Reg2, Reg3 （Reg2とReg3を比較してフラグ更新）
            "101100000001110",  --12: je  14         （一致なら14番地へ）
            "110000000001000",  --13: jmp 8          （無条件で8番地へ戻る）
            "111100000000000",  --14: hlt            （停止）
            "000000000000000"   --15: nop            （何もしない：保険/空き）
        );

begin

    -- ========================================================
    -- PROM読み出し（Fetch段）
    -- ========================================================
    -- CLK_FTの立ち上がりで、PCが指す命令をPROM_OUTへ出す。
    -- ここで出した命令が次のDecode段で解釈されるため、
    -- フェッチ段は “命令ストリームの正しさ” を保証する根幹になる。
    process(CLK_FT)
    begin
        if (CLK_FT'event and CLK_FT = '1') then

            -- ------------------------------------------------
            -- アドレス選択：PC下位4bitでPROMを参照
            -- ------------------------------------------------
            -- MEMが16語なので 0〜15 の範囲に収めるために (3 downto 0) だけ使う。
            -- conv_integer で integer に変換して配列インデックスにする。
            --
            -- 注意：P_COUNTが 0x10,0x20... などでも下位4bitに折り返す。
            PROM_OUT <= MEM(conv_integer(P_COUNT(3 downto 0)));

        end if;
    end process;

end RTL;

-- 【CPU拡張の観点】
-- - 命令数を増やすなら MEMORY のサイズを増やし、P_COUNT全体で参照する。
-- - 分岐やジャンプの正しさを検証するには、PROMに複数パターンのプログラムを入れ替えられる仕組み
--   （別ファイル化/初期化ファイル読み込みなど）があると便利になる。
