-- clk_down.vhd（詳細コメント版）
--
-- 【この回路の目的（CPU設計・FPGA観点）】
-- - 入力クロック CLK_IN を分周して、より遅いクロック CLK_OUT を作る回路である。
-- - FPGAボードの基準クロック（例：50MHz, 100MHz）は人間の目には速すぎるため、
--   自作CPUの bring-up（動作確認）では、
--   - 7セグ表示の変化を目視できる速度に落とす
--   - 命令実行の進み方をゆっくりにしてデバッグしやすくする
--   目的で分周器を噛ませることが多い。
--
-- 【アルゴリズム（分周の本質）】
-- - COUNT を “クロックの立ち上がりごとに 1 ずつ増やす” カウンタとして動かす。
-- - COUNT の各ビットは、入力クロックに対して 2倍・4倍・8倍…と周期が伸びるトグル信号になる。
--
--   たとえば COUNT(0) は毎クロックで 0/1 を反転するので、CLK_IN の 1/2 周波数になる。
--   COUNT(1) は 1/4、COUNT(2) は 1/8 ……
--   つまり COUNT(n) を出力に選ぶと、CLK_IN を 2^(n+1) 分周したクロックが得られる。
--
-- - この設計では COUNT(20) を出力にしているため、分周比は 2^(21) である。
--
-- 【周波数の例（イメージ）】
-- - もし CLK_IN = 50MHz なら、
--     CLK_OUT = 50,000,000 / 2^21 ≒ 23.84 Hz
--   となり、LEDや7セグの更新を目で追えるレベルになる。
--
-- 【CPU設計観点での注意点（重要）】
-- - この方式で作る CLK_OUT は、厳密には “一般的なクロックネットワークに乗った高品質クロック”
--   ではなく、カウンタのビットを直接出しているだけの “分周トグル信号” である。
-- - FPGAでは、クロックはPLL/DCM/Clock Enable で扱うのが推奨であり、
--   ロジックで生成したクロックを別ドメインとして配ると、
--   - スキュー
--   - タイミング制約の難化
--   - 望まないグリッチの扱い
--   などが問題になる場合がある。
--
--   ただし「教育用途」「低速で動かす」「小規模で単純」な自作CPUのデモでは、
--   このような簡易分周器が使われることも多い。
--
-- 【より安全な代替（発展）】
-- - “新しいクロックを作る” のではなく、
--   1) COUNT(20) を Clock Enable（CE）として使い、
--   2) CPUは元のCLK_INで同期しつつ、CE=1の周期だけ状態更新する
--   という方式にすると、クロック品質の問題を避けられる（推奨）。
--
--   ただし、現状の回路は「分周原理の理解」と「目視デバッグ」には十分役立つ。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;  -- COUNT <= COUNT + 1 のために加算演算を許可している（環境によっては非推奨）

-- ============================================================
-- entity：入力クロックを受けて、分周したクロックを出力する
-- ============================================================
entity clk_down is
    port
    (
        CLK_IN  : in  std_logic;  -- 入力クロック（ボードの基準クロック等）
        CLK_OUT : out std_logic   -- 出力クロック（低速化したクロック）
    );
end clk_down;

-- ============================================================
-- architecture：カウンタで分周する
-- ============================================================
architecture RTL of clk_down is

    -- COUNT：分周用カウンタ
    --
    -- 21bit幅（20 downto 0）なので、0〜2^21-1 までカウントしてオーバーフローする。
    -- 各ビットは入力クロックでトグルするため、
    -- COUNT(0) が 1/2、COUNT(1) が 1/4、…、COUNT(20) が 1/2^21 周波数を表す。
    signal COUNT : std_logic_vector(20 downto 0);

begin

    -- --------------------------------------------------------
    -- 分周カウンタの更新（逐次回路）
    -- --------------------------------------------------------
    -- CLK_IN の立ち上がり（'event and = '1'）ごとに COUNT を +1 する。
    -- これにより COUNT は2進カウントアップし、各ビットが規則的に反転する。
    process(CLK_IN)
    begin
        if (CLK_IN'event and CLK_IN = '1') then
            -- 1クロックごとにインクリメント
            -- これが分周の根本：COUNTの上位ビットほどゆっくり反転する
            COUNT <= COUNT + 1;
        end if;
    end process;

    -- --------------------------------------------------------
    -- 分周出力（組合せ代入）
    -- --------------------------------------------------------
    -- COUNT(20) は 2^(20+1)=2^21 分周されたトグル信号。
    -- このビットをそのまま CLK_OUT として外へ出す。
    --
    -- CPUのデモでは、このCLK_OUTをCPUのCLKに入れることで
    -- 命令の進行や表示の更新を遅くして目視確認できる。
    CLK_OUT <= COUNT(20);

end RTL;
