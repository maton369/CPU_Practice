-- d_ff.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 1bitの Dフリップフロップ（D-FF）を記述したものである。
-- - D-FFは「クロック立ち上がり（一般的には）で入力Dを取り込み、出力Qに保持する」記憶素子。
-- - 自作CPUにおいては、D-FFはほぼすべての“状態”の基礎になる。
--   具体例：
--   - レジスタファイル（汎用レジスタ群）
--   - プログラムカウンタ（PC）
--   - 命令レジスタ（IR）
--   - フラグレジスタ（Z/N/C/V等）
--   - パイプラインレジスタ（段間レジスタ）
--   これらは最終的に多数のD-FFの集合として実装される。
--
-- 【回路としての振る舞い（同期回路）】
-- - この回路は組合せ回路ではなく、クロックに同期して状態が更新される「順序回路」である。
-- - クロックの立ち上がりエッジ（rising edge）で、
--     Q_next = D
--   となり、それ以外の時刻では Q は変化しない（保持される）。
--
-- 【VHDLとしてのポイント】
-- - process(CLK) の感度リストに CLK のみを入れることで、
--   クロック変化時のみ評価される“同期プロセス”になる。
-- - `if (CLK'event and CLK = '1') then ...` は
--   「CLKがイベント（変化）した瞬間に、かつ '1' になった時」＝立ち上がり検出。
-- - 近年は `rising_edge(CLK)` の使用が推奨されるが、
--   本コードは古典的な書き方で同じ意味を表している。
--
-- 【自作CPU設計で重要な注意】
-- - D-FFを大量に繋いで“状態”を作ると、クロック境界でデータが確定する。
--   そのためCPUでは「組合せ回路の遅延がクロック周期内に収まるか（タイミング）」が本質になる。
-- - ここでのQ <= D は「非ブロッキング的な信号代入」であり、
--   立ち上がりの瞬間にDをサンプリングし、Qはその後（デルタサイクル）で更新される。
--   これは“同じクロックで複数のレジスタが同時に更新される”というハードウェアの性質に一致する。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic 型を利用するための基本ライブラリ。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity d_ff is
    port
    (
        -- CLK: クロック入力
        -- CPUでは通常、すべての状態要素が同じクロックに同期して更新される。
        CLK : in  std_logic;

        -- D: データ入力（次状態候補）
        -- クロック立ち上がりで取り込まれ、Qに保存される。
        D   : in  std_logic;

        -- Q: データ出力（現在の状態）
        -- クロックが来るまで保持される。
        Q   : out std_logic
    );
end d_ff;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of d_ff is
begin

    -- --------------------------------------------------------
    -- 同期プロセス（クロック立ち上がりで状態更新）
    -- --------------------------------------------------------
    -- 感度リストが CLK のみなので、CLKが変化した時だけプロセスが起動する。
    -- これにより「順序回路（フリップフロップ）」の記述になる。
    process(CLK)
    begin
        -- CLK'event は「CLKに変化があったか」を表す。
        -- かつ CLK='1' のときは、0→1 の立ち上がりエッジである。
        --
        -- 近年の推奨： if rising_edge(CLK) then
        -- だが、意味は同等。
        if (CLK'event and CLK = '1') then

            -- Q <= D は「クロック立ち上がりの瞬間のD」をQに取り込むことを意味する。
            -- 自作CPUの観点では、これが「レジスタに値がラッチされる」動作そのもの。
            --
            -- 重要：
            -- - 信号代入 <= は、同一クロックで複数レジスタが同時更新されるモデルに合う。
            -- - そのため、CPUの状態更新（PC更新、レジスタ書き戻し等）を安全に書ける。
            Q <= D;
        end if;
    end process;

end RTL;

-- 【発展（CPU用レジスタへ）】
-- - 1bit D-FF を N個並べれば Nbitレジスタになる（例：std_logic_vector）。
-- - さらに enable（書き込み許可）や reset（リセット）を追加すると、
--   PC/レジスタ/フラグなど実用的な状態素子になる。
