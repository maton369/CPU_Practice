-- count10_sim.vhd（詳細コメント版：10進カウンタ count10 のテストベンチ）
--
-- 【このファイルの目的（自作CPU観点）】
-- - `count10`（0〜9を繰り返す同期カウンタ）をシミュレーションで検証するテストベンチである。
-- - 自作CPU/SoCでは、カウンタはタイマ・分周・ウェイト生成・表示スキャンなど多用途に使われる。
--   そのため「クロック同期で状態が進む」「リセットで初期状態に戻る」という性質を
--   期待通りに満たすかを、回路単体で確認することが重要である。
--
-- 【テストベンチの検証アルゴリズム（基本形）】
-- 1) DUT（Device Under Test）として count10 を1個インスタンス化する
-- 2) クロック CLK を周期波形として生成する（0/1を交互に繰り返す）
-- 3) リセット RST を所定の時刻でON→OFFして、初期化挙動を確認する
-- 4) 出力 COUNT が
--      - リセット期間中は 0 にクリアされること
--      - リセット解除後に 0→1→…→9→0→… と進むこと
--    を波形で観測する
--
-- 【重要：同期リセットの確認ポイント】
-- - count10 側のRSTは “同期リセット” として実装されている（CLK立ち上がりで評価される）。
-- - したがって、このテストでも
--   「RSTを1にしても、CLK立ち上がりが来るまでCOUNTが変わらない」
--   という挙動が現れるのが正しい。
-- - RSTの波形は 15ns で 1→0 にしているため、
--   ちょうどクロック立ち上がり（例：10ns, 30ns, 50ns...）との関係で
--   “いつリセットが反映されるか” を観測できる。
--
-- 【このTBの刺激設計（時間関係）】
-- - CLKは 20ns周期（10ns Low + 10ns High）を生成している。
--   立ち上がりは 10ns, 30ns, 50ns, ... に発生する。
-- - RSTは
--     t=0〜15ns  : RST=1（リセット要求）
--     t=15ns以降 : RST=0（リセット解除）
--
-- 期待される観測例（同期リセットを前提）：
-- - t=10ns の立ち上がり時点では RST=1 → COUNTは0にクリアされる
-- - t=30ns の立ち上がり時点では RST=0 → COUNTが1に進み始める
--   （初期状態が0で保持されている想定）
--
-- 【注意：このTBのCLK生成プロセスについて】
-- - 現状のCLKプロセスは `process begin ... end process;` の中で
--   0→wait→1→wait の後に末尾へ到達するが、
--   VHDLではプロセスは末尾に到達すると先頭へ戻って繰り返し実行されるため、
--   結果として周期クロックが生成され続ける（よく使う書き方）。
--
-- 【std_logic_unsigned の注意】
-- - TB側では演算をしていないが、教材一式の方針として入っている可能性がある。
-- - 推奨は numeric_std だが、ここでは元コードの方針を踏襲する。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- ============================================================
-- entity: テストベンチは外部ポートを持たない（SIM専用）
-- ============================================================
entity count10_sim is
end count10_sim;

-- ============================================================
-- architecture SIM: シミュレーション用の記述
-- ============================================================
architecture SIM of count10_sim is

    -- --------------------------------------------------------
    -- コンポーネント宣言：DUT（被試験回路）count10
    -- --------------------------------------------------------
    -- 入力：CLK（クロック）, RST（リセット）
    -- 出力：COUNT（0〜9のカウント値）
    component count10
        port
        (
            CLK   : in  std_logic;
            RST   : in  std_logic;
            COUNT : out std_logic_vector(3 downto 0)
        );
    end component;

    -- --------------------------------------------------------
    -- 内部信号：テストベンチ内部の配線
    -- --------------------------------------------------------
    -- CLK/RST は刺激入力（TB側で波形生成する）。
    -- COUNT は観測対象出力（DUTの出力を受ける）。
    signal CLK   : std_logic;
    signal RST   : std_logic;
    signal COUNT : std_logic_vector(3 downto 0);

begin

    -- ========================================================
    -- DUTの実体化（インスタンス化）と配線
    -- ========================================================
    -- count10 を1個置き、TB信号に接続する。
    C1 : count10
        port map(
            CLK   => CLK,
            RST   => RST,
            COUNT => COUNT
        );

    -- ========================================================
    -- クロック生成（stimulus）：CLKの波形
    -- ========================================================
    -- 20ns周期の矩形波を生成する：
    --   0 を 10ns 維持 → 1 を 10ns 維持 → 繰り返し
    --
    -- 自作CPU観点では、ここで作るCLKが “すべての状態更新の基準” になる。
    process
    begin
        CLK <= '0';
        wait for 10 ns;

        CLK <= '1';
        wait for 10 ns;

        -- 末尾に到達するとプロセスは先頭へ戻り、同じ波形を繰り返す。
    end process;

    -- ========================================================
    -- リセット生成（stimulus）：RSTの波形
    -- ========================================================
    -- RST を最初は 1（リセット要求）にし、15ns 後に 0（解除）する。
    -- 同期リセットのため、解除の効果は「次のCLK立ち上がり」から現れるはずである。
    process
    begin
        RST <= '1';         -- リセット要求（初期化したい）
        wait for 15 ns;     -- 15ns 維持

        RST <= '0';         -- リセット解除
        wait;               -- 以降は変化させず停止（観測フェーズ）
    end process;

end SIM;

-- 【テストベンチとしての発展（CPU開発向け）】
-- - COUNTが 0→1→…→9→0 を繰り返すことを assert で自動検証すると回帰試験になる。
-- - リセット解除のタイミングをクロックに揃えたケース/ずらしたケースの両方を試すと、
--   同期リセット設計の意図（クロック境界でのみ初期化される）がより明確に観測できる。
