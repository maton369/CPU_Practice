-- count10.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 0〜9（10進）を繰り返しカウントする 4bit カウンタ（mod-10 counter）である。
-- - CPUコアそのもの（命令実行）ではないが、自作CPU/SoCを作ると必ず出てくる
--   「クロックで進む状態機械（同期回路）」の典型例である。
-- - 具体的な用途例（CPU周辺）：
--   - 7セグ多桁表示のダイナミック点灯（桁選択のスキャン）
--   - タイマ/分周/ウェイト生成（一定回数でイベント発生）
--   - シンプルなステートマシンの周期駆動
--
-- 【アルゴリズム（同期状態更新）】
-- - 立ち上がりクロックごとに COUNT_TMP を次の規則で更新する：
--
--   if RST = 1:
--       COUNT_TMP := 0
--   else if COUNT_TMP = 9:
--       COUNT_TMP := 0
--   else:
--       COUNT_TMP := COUNT_TMP + 1
--
-- - つまり「0→1→2→...→9→0→...」を繰り返す。
-- - これは有限状態機械（FSM）として見ると、状態数10のリング状遷移である。
--
-- 【RSTの扱い（重要）】
-- - 本コードのRSTは “同期リセット” である。
--   理由：
--   - RSTは process(CLK) 内で評価されており、
--     クロック立ち上がりが来たタイミングでのみリセットが反映される。
-- - 非同期リセットにしたい場合は、感度リストに RST を入れたり、
--   if (RST='1') then ... elsif rising_edge(CLK) then ... の形にする必要がある。
--
-- 【std_logic_unsigned の注意】
-- - std_logic_unsigned は std_logic_vector を符号なし整数のように扱って + や比較を可能にする古い拡張。
-- - 近年は numeric_std（unsigned型）を推奨するが、教材ではこの書き方も多い。
-- - 自作CPUで signed/unsigned を明確に扱う段階では numeric_std の方が安全になる。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic / std_logic_vector の基本定義。

use IEEE.std_logic_unsigned.all;
-- std_logic_vector を unsigned とみなして加算（+1）や比較（="1001"）を可能にする拡張。
-- 推奨は numeric_std だが、ここでは元コード方針を踏襲。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity count10 is
    port
    (
        -- CLK: クロック入力
        -- このクロックの立ち上がりごとにカウンタが進む。
        CLK   : in  std_logic;

        -- RST: リセット入力（同期リセット）
        -- RST='1' がクロック立ち上がりでサンプルされるとカウンタを0へ戻す。
        RST   : in  std_logic;

        -- COUNT: 現在のカウント値（4bit）
        -- 0〜9 を表すので4bitで十分。
        -- ただし 10〜15 の値には遷移しない（9の次で0へ戻る）。
        COUNT : out std_logic_vector(3 downto 0)
    );
end count10;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of count10 is

    -- --------------------------------------------------------
    -- 内部信号（状態レジスタ）
    -- --------------------------------------------------------
    -- COUNT_TMP がこの回路の「状態」を保持するレジスタに相当する。
    -- D-FFが4本束ねられた 4bit レジスタ（カウンタレジスタ）と考えられる。
    signal COUNT_TMP : std_logic_vector(3 downto 0);

begin

    -- --------------------------------------------------------
    -- 同期プロセス：クロック立ち上がりで COUNT_TMP を更新
    -- --------------------------------------------------------
    -- 感度リストが CLK のみなので、クロック変化時だけプロセスが起動する。
    -- if (CLK'event and CLK='1') は立ち上がりエッジ検出（rising edge）。
    process(CLK)
    begin
        if (CLK'event and CLK = '1') then

            -- ------------------------------------------------
            -- 1) 同期リセット
            -- ------------------------------------------------
            -- RST='1' のときはカウンタを0に戻す。
            -- ※同期なので、RSTを1にしてもクロックが来るまで反映されない点が重要。
            if (RST = '1') then
                COUNT_TMP <= "0000";

            -- ------------------------------------------------
            -- 2) 9に到達したら0へ戻す（mod-10）
            -- ------------------------------------------------
            -- COUNT_TMP="1001" は 2進数で9。
            -- 0〜9を繰り返すため、9の次のクロックで0に戻す。
            elsif (COUNT_TMP = "1001") then
                COUNT_TMP <= "0000";

            -- ------------------------------------------------
            -- 3) 通常は +1 する
            -- ------------------------------------------------
            -- std_logic_unsigned により COUNT_TMP を unsigned として +1 できる。
            -- 0→1→...→8→9 と進む。
            else
                COUNT_TMP <= COUNT_TMP + 1;
            end if;

        end if;
    end process;

    -- --------------------------------------------------------
    -- 出力への接続
    -- --------------------------------------------------------
    -- COUNT_TMP（内部状態）を外部ポート COUNT に出す。
    -- これにより、外部からは COUNT がカウンタ値として観測できる。
    COUNT <= COUNT_TMP;

end RTL;

-- 【自作CPUでの発展アイデア】
-- - RSTを非同期にしたい場合：プロセスを
--     process(CLK, RST)
--     begin
--       if RST='1' then COUNT_TMP <= "0000";
--       elsif rising_edge(CLK) then ...
--     end
--   のようにする。
-- - さらに enable（カウント許可）を追加すると、タイマ/分周器として使いやすい。
-- - count10 を桁選択に使い、dec_7seg と組み合わせれば多桁7セグ表示の基礎になる。
