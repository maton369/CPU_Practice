maton@Ubuntu22.9530:1770182991