-- and_or.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 1bit入力 A, B に対して AND と OR を同時に出力する組合せ回路である。
-- - 自作CPUでは ALU（算術論理演算器）の一部として、
--   AND/OR のような論理演算は必須級の命令になる。
-- - ここで扱っているのは 1bit だが、CPUでは通常 Nbit（例：16/32bit）なので、
--   この回路をビット幅分だけ並列化（ビットスライス）するか、
--   まとめてベクタ演算（std_logic_vector）に拡張して使うことになる。
--
-- 【VHDLとしてのポイント】
-- - entity: 外部から見える「部品の端子（ポート）」を定義する。
-- - architecture: その部品の「内部動作（回路）」を定義する。
-- - `<=` は信号代入で、ハードウェアの配線関係（同時並行）を表す。
--   ソフトウェアの「順番に実行される代入」とは意味が異なる。
--
-- 【回路としてのポイント】
-- - この記述は完全な組合せ回路（クロック無し）。
-- - 遅延は論理ゲートの伝搬遅延として実装依存で発生する（シミュレーションではデルタサイクル）。
-- - 同時に AND と OR を出しているため、ALU内部で結果候補を並列に作っておき、
--   後段のMUXで命令に応じて選択する設計に繋げやすい。
--
-- 例（ALUの典型構造）：
--   and_result = A AND B
--   or_result  = A OR  B
--   add_result = A + B
--   ...
--   out = MUX(opcode, and_result, or_result, add_result, ...)
--
--   このファイルはその「and_result」「or_result」を作る最小単位の例である。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic / std_logic_vector と、and/or/not などの論理演算子定義を使うために読み込む。
-- 自作CPUでは基本的に std_logic_vector を多用するが、ここでは1bitだけを扱う。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity and_or is
    port
    (
        -- 入力A, B：それぞれ 1bit の論理値
        -- std_logic は '0'/'1' 以外に 'U'(未初期化) や 'Z'(ハイインピーダンス) なども表せる。
        -- 実機回路としては最終的に '0'/'1' に落ちるが、シミュレーションでは未定義状態が見える。
        A      : in  std_logic;
        B      : in  std_logic;

        -- 出力Z_AND：A AND B の結果（1bit）
        Z_AND  : out std_logic;

        -- 出力Z_OR：A OR B の結果（1bit）
        Z_OR   : out std_logic
    );
end and_or;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of and_or is
    -- ここに内部信号（signal）や定数を宣言できる。
    -- 今回は単純な組合せ回路なので内部信号は不要。
begin

    -- --------------------------------------------------------
    -- AND回路
    -- --------------------------------------------------------
    -- `Z_AND <= A and B;`
    --
    -- これは「Z_AND は常に (A AND B) と等しい」という配線を表す。
    -- ソフトウェアのように“この行を実行したら代入が起きる”のではなく、
    -- AやBが変化した瞬間に回路が追従してZ_ANDが変化する（組合せ回路の振る舞い）。
    --
    -- 真理値表（AND）：
    --   A B | Z_AND
    --   0 0 | 0
    --   0 1 | 0
    --   1 0 | 0
    --   1 1 | 1
    Z_AND <= A and B;

    -- --------------------------------------------------------
    -- OR回路
    -- --------------------------------------------------------
    -- `Z_OR <= A or B;`
    --
    -- ORも同様に組合せ回路として常時接続される。
    --
    -- 真理値表（OR）：
    --   A B | Z_OR
    --   0 0 | 0
    --   0 1 | 1
    --   1 0 | 1
    --   1 1 | 1
    Z_OR  <= A or B;

    -- 【自作CPUへの繋げ方（発展）】
    -- - CPUのALUがNbit（例：16bit）なら、A/Bを std_logic_vector(15 downto 0) にして、
    --   `Z_AND <= A and B;` と書くとビットごとのANDが並列に生成される。
    -- - また、AND/ORの結果を直接出すのではなく、
    --   opcodeに応じてどちらかを選ぶMUXを後段に置くのが一般的である。
    --   その場合、このモジュールは「並列に候補を作る部分」として使える。
end RTL;
