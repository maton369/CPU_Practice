-- and_or_sim.vhd（詳細コメント版：テストベンチ / シミュレーション用）
--
-- 【このファイルの目的（自作CPU観点）】
-- - 論理回路 `and_or`（AND/ORゲート）をシミュレーションで検証するための
--   “テストベンチ（testbench）” である。
-- - テストベンチはCPU自作において極めて重要で、
--   ALU・デコーダ・レジスタ・制御回路などを作るたびに、
--   「入力を与えて、出力が期待通りか」を波形で確認する開発ループを支える。
--
-- 【テストベンチのアルゴリズム（考え方）】
-- - DUT（Device Under Test：被試験回路）＝ and_or を1個インスタンス化する
-- - テスト入力（AT, BT）に対して時間変化する波形（刺激 = stimulus）を生成する
-- - DUTの出力（Z_ANDT, Z_ORT）が入力波形に対して正しく反応するかを観測する
--
-- これはCPU開発でも同じで、
--   1) DUT（例：ALU）を置く
--   2) 入力（オペランド、制御信号）を時間で変化させる
--   3) 出力（結果、フラグ）を観測する
-- という検証アルゴリズムが基本になる。
--
-- 【重要：テストベンチは“合成対象ではない”】【SIM専用】
-- - この entity はポートを持たず、外部入出力がない。
-- - wait for 〜 ns といった時間制御はシミュレーション専用で、
--   FPGA合成では通常使えない。
-- - よって architecture 名も SIM としており、明確に“検証用”である。
--
-- 【このテストの波形設計（入力刺激）】
-- - AT は 0 を 10ns 維持 → 1 にして 20ns 維持（その後は指定無し＝プロセス終了）
-- - BT は 0 を 15ns 維持 → 1 にして 20ns 維持（その後は指定無し＝プロセス終了）
--
-- つまり入力の組み合わせは時間によって次のように変化する：
--   t=0〜10ns   : AT=0, BT=0
--   t=10〜15ns  : AT=1, BT=0
--   t=15〜30ns  : AT=1, BT=1
--   t=30〜(終了): 以降はプロセスが止まるので基本的に波形はそのまま保持（ただし観測終了扱いでよい）
--
-- 期待される出力：
-- - Z_ANDT = AT and BT
-- - Z_ORT  = AT or  BT
--
-- 例：
--   (0,0) → AND=0 OR=0
--   (1,0) → AND=0 OR=1
--   (1,1) → AND=1 OR=1


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic を扱うための基本ライブラリ。

-- ============================================================
-- entity: テストベンチは外部ポートを持たない（SIM専用）
-- ============================================================
entity and_or_sim is
end and_or_sim;

-- ============================================================
-- architecture SIM: シミュレーション用の記述
-- ============================================================
architecture SIM of and_or_sim is

    -- --------------------------------------------------------
    -- コンポーネント宣言：DUT（被試験回路）and_or
    -- --------------------------------------------------------
    -- テストベンチ側から見て、and_or は “中身のある回路ブロック”。
    -- これをインスタンス化して入力刺激を与える。
    component and_or
        port
        (
            A     : in  std_logic;
            B     : in  std_logic;
            Z_AND : out std_logic;
            Z_OR  : out std_logic
        );
    end component;

    -- --------------------------------------------------------
    -- 内部信号：テストベンチ内部の配線
    -- --------------------------------------------------------
    -- AT/BT は DUT へ入れる入力信号（刺激波形をここに生成する）。
    -- Z_ANDT/Z_ORT は DUT から出てくる出力信号（観測対象）。
    signal AT     : std_logic;
    signal BT     : std_logic;
    signal Z_ANDT : std_logic;
    signal Z_ORT  : std_logic;

begin

    -- ========================================================
    -- DUTの実体化（インスタンス化）と配線
    -- ========================================================
    -- ここで and_or 回路を 1個置き、テストベンチ信号へ接続する。
    -- 自作CPUの検証でも「DUTを置く→信号を繋ぐ」が常に最初のステップになる。
    C1 : and_or
        port map(
            A     => AT,
            B     => BT,
            Z_AND => Z_ANDT,
            Z_OR  => Z_ORT
        );

    -- ========================================================
    -- 入力刺激（stimulus）生成：AT の波形
    -- ========================================================
    -- process begin ... end process; は無限ループではなく、
    -- この中の記述を上から実行し、wait により時間を進める“シミュレーション専用”の書き方。
    --
    -- ここでは AT を次のように変化させる：
    --   t=0ns   AT=0
    --   t=10ns  AT=1
    --   t=30ns  ここでプロセス終了（以降 AT は 1 のまま）
    process
    begin
        AT <= '0';          -- 初期状態：AT=0
        wait for 10 ns;     -- 10ns 維持
        AT <= '1';          -- AT=1 に切り替え
        wait for 20 ns;     -- 20ns 維持（ここで合計30ns）
        -- ここで process が 끝わるため、以降の刺激は発生しない。
        -- もっと長く試験するなら、最後に wait; を置いて停止させるのが定番。
    end process;

    -- ========================================================
    -- 入力刺激（stimulus）生成：BT の波形
    -- ========================================================
    -- BT を次のように変化させる：
    --   t=0ns   BT=0
    --   t=15ns  BT=1
    --   t=35ns  ここでプロセス終了（以降 BT は 1 のまま）
    process
    begin
        BT <= '0';          -- 初期状態：BT=0
        wait for 15 ns;     -- 15ns 維持
        BT <= '1';          -- BT=1 に切り替え
        wait for 20 ns;     -- 20ns 維持（ここで合計35ns）
        -- 同様に、最後に wait; を置くとシミュレーションを明示的に止められる。
    end process;

end SIM;

-- 【テストベンチとしての発展（CPU設計に近づける）】
-- - 期待値を assert で自動判定すると、波形目視に頼らず回帰試験ができる。
-- - 入力の全組合せ（A,B の 00/01/10/11）を順に流すように波形を設計すると網羅性が上がる。
-- - CPUでは “命令列” をテスト刺激として与え、PC/レジスタ/メモリの期待値を assert で検証する形に拡張できる。
