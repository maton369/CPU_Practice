-- count_nbit.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 任意ビット幅 N_BIT の同期カウンタ（up-counter）である。
-- - クロックの立ち上がりごとに COUNT が +1 され、RST で 0 に戻る。
-- - 自作CPU/SoCでは、可視化・タイマ・分周・待ち状態生成・周期イベント生成など、
--   “一定周期で状態を進める” 機構が頻出であり、汎用Nbitカウンタは周辺回路の基本部品になる。
--
-- 【CPU設計での代表的用途】
-- - タイマ／割り込み源（一定周期で割り込み要求を立てる）
-- - クロック分周（上位ビットを取り出すと遅い周期の矩形波になる）
-- - 7セグ多桁表示のスキャン（桁選択の周期駆動）
-- - デバッグ用“ハートビート”（動作確認の点滅信号）
--
-- 【アルゴリズム（同期状態更新）】
-- - on rising_edge(CLK):
--     if RST = 1:
--         COUNT_TMP := 0
--     else:
--         COUNT_TMP := COUNT_TMP + 1
--
-- - Nbit のため、最大値（2^N - 1）の次は 0 に戻る（自然なオーバーフロー）。
--   これは “mod 2^N カウンタ” であり、CPUではラップアラウンドするカウンタとして扱える。
--
-- 【ジェネリック generic の意味】
-- - VHDLの generic は “パラメータ” に相当する。
-- - N_BIT を変えるだけで、8bitカウンタにも16bitカウンタにもできる。
-- - 自作CPUでは、同じ回路を幅だけ変えて使いたい場面が多く、
--   こうしたパラメタ化は設計資産として強い。
--
-- 【RSTの種類（同期リセット）】
-- - RST は process(CLK) 内で評価されているため同期リセットである。
-- - RST を 1 にしても、クロック立ち上がりが来るまで COUNT_TMP は更新されない。
-- - CPUのリセット戦略（同期/非同期）は全体設計に影響するため、ここは意識点になる。
--
-- 【std_logic_unsigned の注意】
-- - std_logic_unsigned は古い拡張で、std_logic_vector を unsigned とみなして + を可能にする。
-- - 推奨は numeric_std（unsigned型）だが、教材方針としてここでは踏襲している。
-- - CPUで signed/unsigned を厳密に扱う段階では numeric_std 化が望ましい。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity count_nbit is
    generic(
        -- N_BIT: カウンタのビット幅
        -- 既定値は 8（8bitカウンタ）
        -- 例：N_BIT=16 なら 0〜65535 をカウントしてオーバーフローで0に戻る。
        N_BIT : integer := 8
    );
    port(
        -- CLK: クロック入力（立ち上がりで状態更新）
        CLK     : in  std_logic;

        -- RST: リセット入力（同期リセット）
        -- RST='1' がクロック立ち上がりでサンプルされると、カウンタを0に戻す。
        RST     : in  std_logic;

        -- COUNT_N: カウンタ値の出力（N_BIT幅）
        -- LSBが COUNT_N(0)、MSBが COUNT_N(N_BIT-1)。
        COUNT_N : out std_logic_vector(N_BIT - 1 downto 0)
    );
end count_nbit;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of count_nbit is

    -- --------------------------------------------------------
    -- 内部状態レジスタ（カウンタ本体）
    -- --------------------------------------------------------
    -- COUNT_TMP が状態を保持する。
    -- 物理的には N_BIT 本のD-FFで構成されるレジスタの集合と考えられる。
    signal COUNT_TMP : std_logic_vector(N_BIT - 1 downto 0);

begin

    -- --------------------------------------------------------
    -- 同期プロセス：クロック立ち上がりで COUNT_TMP を更新
    -- --------------------------------------------------------
    process(CLK)
    begin
        -- CLK'event and CLK='1' は立ち上がりエッジ検出（rising edge）。
        -- 近年は rising_edge(CLK) を使うことも多いが、意味は同等。
        if (CLK'event and CLK = '1') then

            -- 同期リセット：クロック境界で0に初期化する
            if (RST = '1') then
                -- (others => '0') はベクトル全ビットを0にするVHDLの記法。
                -- N_BITが何であっても一括で0クリアできるので、ジェネリックと相性が良い。
                COUNT_TMP <= (others => '0');

            -- 通常動作：+1 してカウントアップ
            else
                -- N_BIT幅の加算なので、最大値の次はオーバーフローして0へ戻る（mod 2^N）。
                -- 自作CPUで言うと、固定幅レジスタ上の加算と同じ“ラップアラウンド”挙動である。
                COUNT_TMP <= COUNT_TMP + 1;
            end if;

        end if;
    end process;

    -- --------------------------------------------------------
    -- 出力への接続
    -- --------------------------------------------------------
    -- 内部状態（COUNT_TMP）を外部出力（COUNT_N）へ接続する。
    -- デバッグ用途では COUNT_N の特定ビットをLEDに繋ぐと分周器として使える。
    COUNT_N <= COUNT_TMP;

end RTL;

-- 【自作CPUでの発展アイデア】
-- - enable を追加して「カウント停止」「特定条件でのみ+1」を可能にする（タイマ制御に必須）。
-- - terminal count（一定値到達）を検出してパルスを出すと、割り込み源や周期イベントになる。
-- - 上位ビットを取り出すと分周クロックとして使える（例：COUNT_N(N_BIT-1)）。
