-- dec_7seg_sim.vhd（詳細コメント版：7セグデコーダのテストベンチ）
--
-- 【このファイルの目的（自作CPU観点）】
-- - `dec_7seg`（4bit値を7セグ点灯パターンへ変換するデコーダ）を
--   シミュレーションで検証するためのテストベンチ（testbench）である。
-- - 自作CPU開発では「内部の値（レジスタ値/ALU結果/メモリ値）を人間に見える形で出す」
--   ために7セグ表示をよく使う。その際、デコーダが正しく動かないと
--   “CPUが間違っているのか、表示系が間違っているのか” が切り分け不能になる。
-- - したがって、表示系（I/O）の検証を単独で済ませておくことが重要である。
--
-- 【テストベンチの検証アルゴリズム】
-- - DUT（Device Under Test）＝ dec_7seg を1個インスタンス化する
-- - 入力DINを時間経過で 0→1→2→…→15 と順に変化させる（全入力領域の走査）
-- - 出力SEG7が、DINに応じたパターンへ遷移するかを波形で観測する
--
-- 【このTBが“何を網羅しているか”】【網羅性のポイント】
-- - 4bit入力の全組合せ（0〜15）をループで一通り流している。
-- - `dec_7seg` は 0〜9 を数字として定義し、others（10〜15）を全消灯にしている。
--   そのため、このTBでは
--   - 0〜9：定義済みパターンが正しいか
--   - 10〜15：others（全消灯）になっているか
--   の両方を確認できる。
--
-- 【CYCLE（入力更新周期）の意味】
-- - CYCLE = 10ns は「DINを更新する間隔」を表す定数。
-- - テストベンチでは、入力を変える→少し待つ→観測する、という時間刻みを作る必要がある。
-- - dec_7seg は組合せ回路なので理論上は “待たなくても即出力” だが、
--   波形として見やすくするために一定時間維持するのが一般的である。
--
-- 【std_logic_unsigned の注意】
-- - DIN <= DIN + 1 を書くために std_logic_unsigned を使っている。
-- - 近年は numeric_std（unsigned変換）推奨だが、教材方針としてここでは踏襲する。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- ============================================================
-- entity: テストベンチは外部ポートを持たない（SIM専用）
-- ============================================================
entity dec_7seg_sim is
end dec_7seg_sim;

-- ============================================================
-- architecture SIM: シミュレーション用の記述
-- ============================================================
architecture SIM of dec_7seg_sim is

    -- --------------------------------------------------------
    -- コンポーネント宣言：DUT（被試験回路）dec_7seg
    -- --------------------------------------------------------
    -- 4bit入力DINに応じて7bit出力SEG7を生成するデコーダ。
    component dec_7seg
        port
        (
            DIN  : in  std_logic_vector(3 downto 0);
            SEG7 : out std_logic_vector(6 downto 0)
        );
    end component;

    -- --------------------------------------------------------
    -- 定数：入力を更新する周期（シミュレーションの時間刻み）
    -- --------------------------------------------------------
    -- 10nsごとにDINを更新し、波形上で各入力値が一定時間保持されるようにする。
    constant CYCLE : time := 10 ns;

    -- --------------------------------------------------------
    -- 内部信号：テストベンチ内部の配線
    -- --------------------------------------------------------
    -- DIN は刺激入力。初期値 "0000"（0）から開始する。
    -- SEG7 は観測対象出力。
    signal DIN  : std_logic_vector(3 downto 0) := "0000";
    signal SEG7 : std_logic_vector(6 downto 0);

begin

    -- ========================================================
    -- DUTの実体化（インスタンス化）と配線
    -- ========================================================
    -- dec_7seg を1個置き、TB内部信号へ接続する。
    C1 : dec_7seg
        port map(
            DIN  => DIN,
            SEG7 => SEG7
        );

    -- ========================================================
    -- 入力刺激（stimulus）生成：DIN を 0〜15 まで順に変化
    -- ========================================================
    -- このプロセスはシミュレーション専用の時間制御を行う。
    --
    -- for I in 0 to 15 loop
    --   wait for CYCLE;   （一定時間その値を保持）
    --   DIN <= DIN + 1;   （次の値へインクリメント）
    -- end loop;
    --
    -- これによりDINは
    --   0,1,2,...,15
    -- と全パターンを一通り通過する（網羅試験になっている）。
    process
    begin
        -- I はループ回数のための変数であり、DIN自体は DIN<=DIN+1 で更新している。
        -- ここでは “入力空間を走査する” というテストベンチの典型形になっている。
        for I in 0 to 15 loop
            wait for CYCLE;     -- 現在のDINを一定時間保持して観測可能にする
            DIN <= DIN + 1;     -- 次の入力値へ進める（4bitなので 15+1=0 に戻るが、loopはここで終了）
        end loop;

        -- wait; は無期限待機（これ以上刺激を出さず、シミュレーションをここで止める）に相当する。
        -- ツール上ではこの時点で波形を見て結果確認できる。
        wait;
    end process;

end SIM;

-- 【テストベンチとしての発展（CPU開発向け）】
-- - 目視だけでなく assert を入れると自動判定でき、回帰試験に強くなる。
--   例：DIN="0011" のとき SEG7 が "0110000" か、などを時刻ごとにチェックする。
-- - 7セグの“ビット並び/極性”はボード依存なので、実機に合わせた期待値表を
--   テストベンチ側にも持たせると、表示系の不一致を早期に検出できる。
