-- half_adder.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 1bit入力 A, B の「足し算」を行い、
--     S  : Sum（和の下位1bit）
--     CO : Carry Out（桁上がり）
--   を出力する「半加算器（Half Adder）」である。
--
-- - 自作CPUのALU（算術論理演算器）では加算（ADD）が最重要命令の1つであり、
--   Nbit加算器（例：16/32bit）の基本部品として半加算器/全加算器は頻出である。
-- - 半加算器は「Carry In（入力桁上がり）」を扱わない加算器なので、
--   多ビット加算器を作るには通常「全加算器（Full Adder）」を連結する。
--   ただし、最下位ビット（LSB）は Carry In = 0 なので、LSBだけ半加算器で始める設計もできる。
--
-- 【VHDLとしてのポイント】
-- - entity: 外部インタフェース（ポート：端子）の宣言
-- - architecture: 内部回路（論理式・配線）の記述
-- - `<=` は信号代入で、ソフトウェアの逐次実行ではなく「回路の接続（同時並行）」を表す。
--
-- 【半加算器の論理】
-- - 1bitの加算は次の真理値表で表される。
--
--   A B | S CO
--   ----+------
--   0 0 | 0  0
--   0 1 | 1  0
--   1 0 | 1  0
--   1 1 | 0  1
--
-- - ここから論理式は次のように導ける。
--   - S  = A ⊕ B   （xor：排他的論理和）
--   - CO = A ∧ B   （and：両方1のときだけ桁上がり）
--
-- 【CPU設計への接続（発展）】
-- - Nbit加算器：
--   - LSBは half_adder（Carry In = 0）でも良い
--   - それ以外は full_adder（Carry In を考慮）を連結するのが一般的
-- - ALUでは、加算結果だけでなくフラグ（Z/N/C/Vなど）も必要になるので、
--   CO（キャリ）や最上位ビットの変化を使ってフラグ生成へ繋げる。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic 型と、and/xor などの論理演算子を利用するために読み込む。
-- CPU回路では std_logic_vector（多ビット）へ拡張するのが一般的。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity half_adder is
    port
    (
        -- 入力A, B：1bit
        -- std_logic は 0/1 以外も表せる（U, X, Z等）。
        -- シミュレーションで未初期化を検出できるので、CPUの回路検証で役に立つ。
        A  : in  std_logic;
        B  : in  std_logic;

        -- 出力S：和（Sum）
        -- 1bit加算の「下位bit」に相当する。
        S  : out std_logic;

        -- 出力CO：Carry Out（桁上がり）
        -- A=B=1 のときに 1 になる。
        -- 多ビット加算器では、このCOが次段のCarry Inに接続される。
        CO : out std_logic
    );
end half_adder;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of half_adder is
    -- 内部信号が必要ならここで宣言できるが、今回は不要（論理式が直接書ける）。
begin

    -- --------------------------------------------------------
    -- S（Sum）の生成
    -- --------------------------------------------------------
    -- S <= A xor B;
    --
    -- 排他的論理和（XOR）は
    -- - AとBが異なるときに1
    -- - AとBが同じときに0
    -- となるため、1bit加算の「下位bit」と一致する。
    --
    -- 自作CPU観点：
    -- - 加算器内部でXORは非常によく使われる。
    -- - XORゲートの実装コストや遅延は、加算器の速度（クリティカルパス）に影響する。
    S <= A xor B;

    -- --------------------------------------------------------
    -- CO（Carry Out）の生成
    -- --------------------------------------------------------
    -- CO <= A and B;
    --
    -- ANDは A=B=1 のときだけ1になるため、
    -- 1bit加算で桁上がりが発生する条件（1+1=10）と一致する。
    --
    -- 自作CPU観点：
    -- - Carryは多ビット加算器の連鎖に関わり、速度のボトルネックになりやすい。
    -- - 高速化したい場合、リップルキャリーではなく
    --   キャリー先読み（Carry Lookahead）等の構造へ発展する。
    CO <= A and B;

end RTL;
