-- clk_gen.vhd（詳細コメント版：ステージクロック生成 / 段階実行のタイミング制御）
--
-- 【このモジュールの目的（CPU設計観点）】
-- - ベースクロック `CLK` を入力として、
--   CPUの各ステージ（Fetch / Decode / Execute / WriteBack）を順番に動かすための
--   “ワンホット（one-hot）なステージクロック” を生成する。
--
-- - 具体的には、ベースクロックの立ち上がりごとに
--   CLK_FT → CLK_DC → CLK_EX → CLK_WB →（再び）CLK_FT …
--   の順で「どれか1本だけが '1' になる」ように出力を切り替える。
--
-- 【この方式の意味（段階実行のアルゴリズム）】
-- - 通常のパイプラインCPUは、全ステージが同一クロックで並列に動く（各段が同時に更新）ことが多い。
-- - 一方この設計は「1クロックごとに実行段を切り替える」方式で、
--   1命令を 4 サブサイクル（FT/DC/EX/WB）に分けて逐次的に進めるイメージになる。
--
--   段階実行の1命令（概念）：
--   - FT: 命令をROMから読む
--   - DC: 命令をデコードし、レジスタ/RAMの読み出し準備
--   - EX: ALU/分岐/ロードストア制御を実行し、書き戻しデータを生成
--   - WB: レジスタ/RAMへ書き戻し
--
-- - 自作CPUでは、まずこのように“逐次で確実に動く”設計にすると
--   タイミングの難易度を下げられ、デバッグもしやすい。
--
-- 【重要：これは「クロックゲーティング」に近い】
-- - 出力は “CLKの分周クロック” ではなく、「ステージイネーブル（enable）」として使うのが本質。
-- - FPGA/ASIC設計の一般論では、クロックを論理で直接ON/OFFするのは注意が必要で、
--   可能なら “同一クロック + enable” にするのが安全である。
-- - ただし教材/小規模CPUでは、段のトリガとして擬似クロックを配る設計が採られることがある。
--   この場合、配線遅延やグリッチが起きないように
--   「完全に同期的に '0'/'1' を切り替えているか」が重要になる。
--
-- 【この回路の生成アルゴリズム（実装の中身）】
-- - 2bitカウンタ COUNT を持ち、CLK立ち上がりごとに +1 する。
-- - COUNT の値で case 分岐し、対応する出力だけ '1'、残りを '0' にする。
--
--   COUNT="00" → FT=1
--   COUNT="01" → DC=1
--   COUNT="10" → EX=1
--   COUNT="11" → WB=1
--
-- - これにより、4段のワンホットシーケンスが完成する。
--
-- 【観測上の注意（波形としてどう見えるか）】
-- - 各出力は “1ベースクロック周期だけ '1' になるパルス” のように見える。
-- - つまり、FT/DC/EX/WB はそれぞれベースクロックの1/4周期で“有効化”される。
-- - CPU全体では、1命令を完了するのにベースクロック4サイクル相当がかかる設計になる。
--
-- 【リセットが無い点の注意】
-- - COUNT の初期値は "00" に初期化されているため、シミュレーション上は
--   最初の立ち上がりで FT が '1' から始まる。
-- - 実機（FPGA）では初期値が確実に入るかはデバイス/合成設定に依存する場合がある。
--   堅牢にするなら RESET_N などで COUNT と出力を既知状態へ初期化するのが定石である。


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- ============================================================
-- entity: ベースクロック → ステージクロック（ワンホット）生成
-- ============================================================
entity clk_gen is
    port
    (
        CLK     : in  std_logic;  -- ベースクロック
        CLK_FT  : out std_logic;  -- Fetch段を動かすトリガ
        CLK_DC  : out std_logic;  -- Decode段を動かすトリガ
        CLK_EX  : out std_logic;  -- Execute段を動かすトリガ
        CLK_WB  : out std_logic   -- WriteBack段を動かすトリガ
    );
end clk_gen;

-- ============================================================
-- architecture RTL: 2bitカウンタで4段を順番に有効化
-- ============================================================
architecture RTL of clk_gen is

    -- --------------------------------------------------------
    -- COUNT: 2bitの段カウンタ
    -- --------------------------------------------------------
    -- "00"→"01"→"10"→"11"→"00"... と循環し、
    -- その値に応じて出力のワンホットパターンを切り替える。
    signal COUNT : std_logic_vector(1 downto 0) := "00";

begin

    -- ========================================================
    -- CLK立ち上がりで段を進める順序回路
    -- ========================================================
    process(CLK)
    begin
        -- 立ち上がりエッジ検出（同期回路の基本形）
        if (CLK'event and CLK = '1') then

            -- ------------------------------------------------
            -- 現在のCOUNTに応じて、どの段を有効化するかを決定
            -- ------------------------------------------------
            -- ここでは “必ず1本だけ '1'” になるようにしている。
            case COUNT is

                -- Fetch段だけ有効
                when "00" =>
                    CLK_FT <= '1';
                    CLK_DC <= '0';
                    CLK_EX <= '0';
                    CLK_WB <= '0';

                -- Decode段だけ有効
                when "01" =>
                    CLK_FT <= '0';
                    CLK_DC <= '1';
                    CLK_EX <= '0';
                    CLK_WB <= '0';

                -- Execute段だけ有効
                when "10" =>
                    CLK_FT <= '0';
                    CLK_DC <= '0';
                    CLK_EX <= '1';
                    CLK_WB <= '0';

                -- WriteBack段だけ有効
                when "11" =>
                    CLK_FT <= '0';
                    CLK_DC <= '0';
                    CLK_EX <= '0';
                    CLK_WB <= '1';

                -- 想定外の値（基本的に起きないが保険）
                when others =>
                    null;
            end case;

            -- ------------------------------------------------
            -- 次の段へ進める（2bitなので4周期で一周する）
            -- ------------------------------------------------
            COUNT <= COUNT + 1;

        end if;
    end process;

end RTL;

-- 【CPU設計としての次の検討ポイント】
-- - RESET_N を追加して、COUNTと出力を確実に既知状態へ初期化する（実機で強い）。
-- - 出力を “クロック” として扱うより “enable” として扱う設計に寄せると安全性が上がる。
--   （同一CLKで全段を駆動し、段ごとに enable で更新する方式）
