-- adder_4bit_lib.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 4bit入力 AIN, BIN を加算し、5bit出力 SOUT に結果を出す加算器である。
-- - ただし、前回の adder_4bit.vhd のように half_adder / full_adder を接続して
--   “構造として加算器を作る” のではなく、
--   VHDLの演算子「+」を使って “振る舞い（behavior）として加算” を記述している。
--
-- - 自作CPUを作る観点では、これは次の違いとして重要である。
--   1) 構造記述（ゲート/加算器セルを繋ぐ）：
--      - キャリー鎖や遅延が見えやすい
--      - ハードウェアの作りを学ぶのに向く
--   2) 振る舞い記述（+ 演算子で書く）：
--      - 設計が短く、可読性が高い
--      - 合成ツールが内部で最適な加算器（キャリー鎖/専用キャリーチェーン等）を生成する
--      - “自作CPUのALUを作る” という目的では実務的にこちらが多い
--
-- 【重要：std_logic_unsigned の意味と注意】
-- - std_logic_unsigned は「std_logic_vector を符号なし整数として扱い、+ などを使えるようにする」
--   ための古い拡張ライブラリである。
-- - 近年の推奨は IEEE.numeric_std を使い、
--   unsigned/signed 型に明示変換する書き方である（移植性と明確さが上がる）。
-- - ただし教材としては std_logic_unsigned を使う例も多いので、
--   ここでは原文を尊重して維持しつつ、意味をコメントで明示する。
--
-- 【なぜ出力が5bitなのか】
-- - 4bitの最大値は 15（1111）
-- - 15 + 15 = 30（11110）なので、結果は最大で5bit必要。
-- - そのため、入力の前に '0' を連結して 5bit化してから加算している。
--   これは「桁あふれ（キャリーアウト）を結果に含める」ための典型手法である。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic / std_logic_vector の定義と論理演算子を使うために読み込む。

use IEEE.std_logic_unsigned.all;
-- std_logic_vector を “符号なし（unsigned）” とみなして + などの算術演算を許可する拡張。
-- 注意：現在は numeric_std（unsigned型）を推奨することが多い。
--       ただし、このファイルは “短く加算を書く” ことを目的にこのライブラリを使用している。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity adder_4bit_lib is
    port(
        -- 4bit入力（LSBが(0), MSBが(3)）
        AIN  : in  std_logic_vector(3 downto 0);
        BIN  : in  std_logic_vector(3 downto 0);

        -- 5bit出力（桁あふれを含む）
        -- SOUT(3 downto 0) が和の下位4bit、
        -- SOUT(4) が最上位キャリー（桁あふれ）に相当する。
        SOUT : out std_logic_vector(4 downto 0)
    );
end adder_4bit_lib;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of adder_4bit_lib is
begin

    -- --------------------------------------------------------
    -- 5bit化して加算する（桁あふれを保持するため）
    -- --------------------------------------------------------
    -- SOUT <= ('0' & AIN) + ('0' & BIN);
    --
    -- ('0' & AIN) は 1bit '0' を上位側に付け足して 5bit に拡張する操作。
    -- 例：AIN="1010"(10) → ('0' & AIN)="01010"(10)
    --
    -- これを両入力に対して行うことで、
    -- 4bit同士の加算で生じる「最上位のキャリー」を結果のbit4に保持できる。
    --
    -- 自作CPU観点：
    -- - これは ALU の Carry Flag（Cフラグ）に相当する情報を出力に含める操作と考えられる。
    -- - 構造記述（full_adder連結）では CO がチェーンの最後に出てくるが、
    --   振る舞い記述ではこのようにビット幅を増やすことでキャリーを“見える化”できる。
    --
    -- 合成（FPGA/ASIC）では、ツールが内部で加算器回路を生成する。
    -- FPGAなら専用のキャリーチェーン資源が使われ、高速な実装になりやすい。
    SOUT <= ('0' & AIN) + ('0' & BIN);

end RTL;

-- 【参考：より推奨される numeric_std 版の考え方（説明のみ）】
-- - numeric_std を使う場合は、
--     unsigned('0' & AIN) + unsigned('0' & BIN)
--   のように型を明示し、結果を std_logic_vector に戻すのが定石である。
-- - “CPUを作る” という観点では、符号付き/符号なしを明確に区別できるため、
--   特にSUBや比較、オーバーフロー判定を扱う段階で numeric_std の方が安全になる。
