-- dec_7seg.vhd（詳細コメント版）
--
-- 【このモジュールの目的（自作CPU観点）】
-- - 4bit入力（DIN）を、7セグメントLED表示用の7bit信号（SEG7）へ変換するデコーダである。
-- - 自作CPUを作るとき、演算結果やレジスタ値を「人間が見える形」に出す仕組みが必要になる。
--   その最小で分かりやすい出力デバイスが 7セグ表示であり、
--   この回路は「数値(0〜9) → セグ点灯パターン」への変換を担当する。
--
-- 【CPU設計での位置づけ】
-- - CPUコア（ALU/レジスタ/制御）そのものではなく、“I/O周辺回路” に相当する。
-- - ただし bring-up（初期動作確認）では、
--   - メモリの特定アドレスに書いた値を表示する
--   - レジスタの値を表示する
--   といった用途で非常に役立つため、デバッグ用の観測点として重要である。
--
-- 【7セグメントの基本】
-- - 7セグは通常 a,b,c,d,e,f,g の7本のLEDセグメントで数字を表す。
-- - `SEG7` は 7bit（6 downto 0）で、どのビットがどのセグメントに対応するかは
--   ボード配線（制約ファイル）によって決まる。
-- - さらに、7セグには
--   - 共通アノード（Common Anode）
--   - 共通カソード（Common Cathode）
--   の2種類があり、「0で点灯 / 1で点灯」が逆になる。
-- - このコードでは "0" が点灯、"1" が消灯になっているパターンが多いので、
--   一般的には “アクティブLow（0で点灯）” の配線を想定していると考えられる。
--   （ただし最終的にはボード仕様に合わせてビット並びと極性を確認する必要がある）
--
-- 【回路としての性質】
-- - process(DIN) の感度リストに DIN が入っているため、
--   DIN が変化するたびに case 文が評価される。
-- - これは「組合せ回路（コンビ回路）」としてのデコーダであり、
--   クロックや状態（レジスタ）を持たない。
-- - 言い換えると、DIN を入力した瞬間に対応するセグパターンが出力される（遅延は実装依存）。
--
-- 【対応範囲】
-- - "0000"〜"1001"（0〜9）を表示対象としている。
-- - それ以外（10〜15）は others で "1111111"（全消灯）としている。
--   bring-up用途では “未定義値を表示しない/誤解させない” という意味で妥当である。


library IEEE;
use IEEE.std_logic_1164.all;
-- std_logic / std_logic_vector を扱うための基本ライブラリ。

-- ============================================================
-- entity: 入出力（ポート）の宣言
-- ============================================================
entity dec_7seg is
    port
    (
        -- 4bit入力：表示したい値（0〜15の範囲を取り得る）
        -- 自作CPUでは「レジスタ値の下位4bit」や「I/Oに書いた値」をここに入れる想定。
        DIN  : in  std_logic_vector(3 downto 0);

        -- 7bit出力：7セグ表示の点灯パターン
        -- どのビットが a〜g のどれに対応するかはボード配線に依存。
        -- また、0で点灯（active-low）か1で点灯（active-high）かも配線に依存。
        SEG7 : out std_logic_vector(6 downto 0)
    );
end dec_7seg;

-- ============================================================
-- architecture: 回路（内部実装）の記述
-- ============================================================
architecture RTL of dec_7seg is
begin

    -- --------------------------------------------------------
    -- 組合せデコーダ（DIN → SEG7）
    -- --------------------------------------------------------
    -- process(DIN) としているので、DIN が変化するたびに内部が再評価される。
    -- クロックが無いので“同期回路”ではなく“組合せ回路”になる。
    process(DIN)
    begin
        -- case 文で DIN の値ごとに対応する7セグパターンを割り当てる。
        --
        -- 各パターン文字列（例："1000000"）の意味：
        -- - 7本のセグメントそれぞれを点灯/消灯させるビット列。
        -- - この例は多くの場合 active-low（0で点灯）を想定した表現になっている。
        --
        -- 注意：
        -- - 実際にどのセグが点灯するかは “ビット順序（SEG7(6)がaなのかgなのか等）” に依存する。
        -- - ここでは「このボード配線で数字が正しく見える」ように既に決め打ちされた表だと解釈する。
        case DIN is
            -- 0 を表示（通常は a,b,c,d,e,f 点灯 / g 消灯）
            when "0000" => SEG7 <= "1000000";

            -- 1 を表示（通常は b,c 点灯）
            when "0001" => SEG7 <= "1111001";

            -- 2 を表示
            when "0010" => SEG7 <= "0100100";

            -- 3 を表示
            when "0011" => SEG7 <= "0110000";

            -- 4 を表示
            when "0100" => SEG7 <= "0011001";

            -- 5 を表示
            when "0101" => SEG7 <= "0010010";

            -- 6 を表示
            when "0110" => SEG7 <= "0000010";

            -- 7 を表示
            when "0111" => SEG7 <= "1111000";

            -- 8 を表示（通常は全点灯）
            when "1000" => SEG7 <= "0000000";

            -- 9 を表示
            when "1001" => SEG7 <= "0010000";

            -- 10〜15（A〜F相当）や不定値は表示しない（全消灯）：
            -- bring-upでは「想定外の値を出さない」方がバグの切り分けがしやすいことが多い。
            when others => SEG7 <= "1111111";
        end case;
    end process;

end RTL;

-- 【自作CPUでの実用上の発展】
-- - 7セグが複数桁ある場合は、各桁を高速に切り替える “ダイナミック点灯（多重化）” が必要。
--   その場合は、
--   - 表示したい多ビット値を各4bit（ニブル）に分解
--   - dec_7seg を桁ごとに使う（または共有してMUX）
--   - 桁選択信号をタイマで回す
--   という構造になる。
-- - CPUのデバッグ用途なら「PC」「IR」「レジスタ」などを切り替え表示できるようにすると強い。
